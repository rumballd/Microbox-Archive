--
-- MON09 monitor ROM for the MB2K 
-- Version 1.0	 31-3-05	   (6Kbyte ROM using three block RAMs)
--
library IEEE, UNISIM;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use UNISIM.vcomponents.all;
		
entity MON09_rom is
    Port (
       clk   : in  std_logic;
	  rst   : in  std_logic;
	  cs    : in  std_logic;
	  rw    : in  std_logic;
       addr  : in  std_logic_vector (12 downto 0);
       rdata : out std_logic_vector (7 downto 0);
       wdata : in  std_logic_vector (7 downto 0)
    );
end MON09_rom;
 
architecture Behavioral of MON09_rom is

   -- RAMB16_S9: Virtex-II/II-Pro, Spartan-3 2k x 8 + 1 Parity bit Single-Port RAM
   -- Xilinx  HDL Language Template version 6.3.1i

   signal dp0, dp1, dp2 : std_logic_vector(0 downto 0);	-- loop parity bit output to input
   signal we, cs0, cs1, cs2 : std_logic;
   signal rdata0, rdata1, rdata2 : std_logic_vector(7 downto 0);

begin
   
   RAM_0 : RAMB16_S9    -- $E800 - EFFF
   generic map (
      INIT => X"000", --  Value of output RAM registers at startup
      SRVAL => X"000", --  Ouput value upon SSR assertion
      WRITE_MODE => "WRITE_FIRST", --  WRITE_FIRST, READ_FIRST or NO_CHANGE
    INIT_00 => x"3595AD588CDFF630E88EFC27EC8D1434963595AD83E8BD588CDFF63CE88E1634",
    INIT_01 => x"83E87DE872E867E863E858E84DE842E8943595AD588DDFF636E88E1434ED8D94",
    INIT_02 => x"B6EE270185E0E7B639A1E7B6F9270185A0E7B63991E7B6F927018590E7B689E8",
    INIT_03 => x"90E7B639A1E7B7EE2702C5E0E7F639A1E7B7F92702C5A0E7F6397C001739A1E7",
    INIT_04 => x"D4E7B7D3E7B7D2E7B74FD1E7B703861634390184E0E7B6390184A0E7B6390184",
    INIT_05 => x"7FB8DF7F9635D3E77FD2E77FC7DF7FB7DF7FB8DF7FF62618C15C168DD3E7F75F",
    INIT_06 => x"F22650C15CD0E7B7B8DFF7D2E7F72086B8DFF6063439D2E77FB8DF7F078DD2E7",
    INIT_07 => x"F703C60520D1E7F730C607278085252520812720B7E9BD0527C7DF7D76348635",
    INIT_08 => x"B696AD482FE98E1634F635D2E7B7B8DFB7062750814CB8DFB6D0E7B77F84D1E7",
    INIT_09 => x"E93EF49DE99DE99DE99DE99DE99DE99DE9E6201635D3E7B7B7DFB6D2E7B7B8DF",
    INIT_0a => x"E9E5E9DFE99DE99DE99DE99DE99DE99DE9B0E9B7E9B3E98FE89EE985E979E96F",
    INIT_0b => x"2750814CB8DFB639B8DFB7032B4AB8DFB69DE99DE99DE99DE99DE9BCE8CBE89D",
    INIT_0c => x"DFB639B7DFB7BCE87ED3E7B7B7DFB717865C8D0D2618814CB7DFB639B8DFB703",
    INIT_0d => x"F702C606265DC7DFF639B8DF7FB7DF7FBCE87ED3E7B7B7DFB74F528DF62A4AB7",
    INIT_0e => x"8639C7DF7AD2E7B7B8DFB7208039C7DF7AD3E7B7B7DFB720800C2602C139C7DF",
    INIT_0f => x"1786022A4AD4E7B639D4E7B74F012618814CD4E7B639D1E7B7038639D1E7B730",
    INIT_10 => x"2BEB2BEBF4EAE8EA54EA54EA54EAA4EAA4EAA4EAA4EAA4EABEEA5FEA39D4E7B7",
    INIT_11 => x"54EA54EA54EA54EA54EA54EA54EA54EA54EA54EA54EA54EA54EA2BEB2BEB2BEB",
    INIT_12 => x"3439011A5D40C639FE1C5D5F54EA54EA54EA28EC28EC28EC28EC23ECC3EB54EB",
    INIT_13 => x"C0E7B74FF9265AA0A780A65F80DE8E1000008EC1E7F7C0E7B7028B318D103420",
    INIT_14 => x"0435011F3D0AC604345ABEFF162035F9265A80A7A0A65F80DE8E101035C1E7B7",
    INIT_15 => x"023439011A5D80C69CFF16032655AA831080DEFCB38D80DE8E01C64F39101F3A",
    INIT_16 => x"0635F9265AA0A780A65F80DE8E1006342034023559EA7E02350526408480E7B6",
    INIT_17 => x"A780A65F80DE8E100634203473FF16048B57001710342034220016028BB3FF17",
    INIT_18 => x"4FF9265A80A7A0A65F80DE8E1000008EC1E7F7C0E7B7048B3E8D0635F9265AA0",
    INIT_19 => x"14FF16032655AA831080DEFCB4FF1780DE8E01C64F29FF162035C1E7B7C0E7B7",
    INIT_1a => x"7386CCDF7FCBDF7F0234043439101F3A0435011F3D24C604345A39011A5D80C6",
    INIT_1b => x"2441ECBD5F36245FECBD02353D245FECBD023544245FECBD8EDFB64C245FECBD",
    INIT_1c => x"35891F142441ECBD02341B2441ECBDEB265ACBDF7C0324CCDFB7CCDFBB80A730",
    INIT_1d => x"DFF709C6F5245FECBD1586092010C60D205F03245FECBD06860E26CBDFB31002",
    INIT_1e => x"ECBD0235D5245FECBD8EDFB6DD245FECBD7286CCDF7FCBDF7F02340434395DCB",
    INIT_1f => x"EB265ACBDF7C0324CCDFB7CCDFBBBF245FECBD80A65FC7245FECBD0235CE245F",
    INIT_20 => x"DFF70AC602205F032606819C2441ECBDA1245FECBDCCDFB6A9245FECBDCBDFB6",
    INIT_21 => x"5D011A10C604205F03260681072441ECBD0C245FECBD5186395DCBDFF6395DCB",
    INIT_22 => x"34B035A1E7B6B035EE261F30F6263F310A2547A0E7B6E2048E10E8038E303439",
    INIT_23 => x"B70235B0350235ED261F30F5263F310C254747A0E7B6E2048E10E8038E023430",
    INIT_24 => x"8EDFF703E63034A7DF9F6E390127078DA5DF9F6EA3DF9F6EA1DF9F6EB035A1E7",
    INIT_25 => x"A614C6A1DF8E108B3004EA8E3D14C639011A5D0FC630350826FF8185A69DDF8E",
    INIT_26 => x"AD0425BC8D8BDF8E8EDFB74FADDF9F6EABDF9F6EA9DF9F6E3035F9265AA0A780",
    INIT_27 => x"2C8D80E7B7038A80E7B60234B3DF9F6EB1DF9F6E39EA2604814C8EDFB6AFDF9F",
    INIT_28 => x"E7B7028A108D80E7B7FE8480E7B6023482351E8D80E7B7FD84258D80E7B7FE84",
    INIT_29 => x"008E80E7F61434B635FB263F313D29008E1036348235028D80E7B7018A098D80",
    INIT_2a => x"261F30CF8D80E7F7FDC4D68D80E7F702CADD8D80E7F701CA0220FEC404254808",
    INIT_2b => x"01C480E7F6B18D80E7F703CA4808008E4FBD8D80E7F701CA80E7F614349435E0",
    INIT_2c => x"80E7F701CA80E7F604349435DF261F309C8D80E7F7FDC401CA80E7F6018A0227",
    INIT_2d => x"1780E7F701CA80E7F60434843579FF1780E7F7FDC481FF1780E7F702CA89FF17",
    INIT_2e => x"00000000000000000000000084355AFF1780E7F7FDC462FF1780E7F702CA6AFF",
    INIT_2f => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_30 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_31 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_32 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_33 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_34 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_35 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_36 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_37 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_38 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_39 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3a => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3b => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3c => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3d => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3e => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3f => x"0000000000000000000000000000000000000000000000000000000000000000"



	 )

   port map (
      DO => rdata0,                -- 8-bit Data Output
      DOP => dp0,                  -- 1-bit parity Output
      ADDR => addr(10 downto 0),   -- 11-bit Address Input
      CLK => clk,                  -- Clock
      DI => wdata,                 -- 8-bit Data Input
      DIP => dp0,                  -- 1-bit parity Input
      EN => cs0,                   -- RAM Enable Input
      SSR => rst,                  -- Synchronous Set/Reset Input
      WE => we                     -- Write Enable Input
   );
   -- End of RAMB16_S9_inst instantiation
   
   RAM_1 : RAMB16_S9    -- $F000 - $F7FF
   generic map (
      INIT => X"000", --  Value of output RAM registers at startup
      SRVAL => X"000", --  Ouput value upon SSR assertion
      WRITE_MODE => "WRITE_FIRST", --  WRITE_FIRST, READ_FIRST or NO_CHANGE
    INIT_00 => x"87F37DF35EF339F32EF31DF369F200F3EDF2F9F223E800E821E810E82CF2A4F0",
    INIT_01 => x"ECECD4ECD0ECCCEC99EC90EC8CEC88EC84EC11F305F38EF389F34BF34FF385F3",
    INIT_02 => x"69F269F269F269F269F269F269F269F269F269F23EF41DF4F1F319F4EDF3F0EC",
    INIT_03 => x"42E869F269F269F269F269F269F269F269F269F269F269F269F269F269F269F2",
    INIT_04 => x"B5ED96ED63ED39ED10EDF4ECD5F3BCF3B1F369F269F269F269F269F269F269F2",
    INIT_05 => x"106FDECE109CDFB7AA86F92600E08C80A780DF8E4F1027AA819CDFB641EC5FEC",
    INIT_06 => x"F2BE80E7B70386C1E7B7C0E7B74FF8268CDF8C80AF1082DF8E5EF28E1080DFFF",
    INIT_07 => x"BD0EC6B5DF7F8DDFF701C454891F8CDFF701C4891F4444444480E7B698DFBF34",
    INIT_08 => x"8D0016B5DFB7FF860827AA81F1F3BD0EC61DF4BD0EC6AA86A5002710AA81F1F3",
    INIT_09 => x"076E20B5DF7FF62640C15C1DF4BD80A65F6EF18E1DF3BDB80B8E00F3BD3FF18E",
    INIT_0a => x"6964616F6C6572202C435452206E69206572756C696166207265776F50070707",
    INIT_0b => x"010077AA0000000000000005013102090000040D0A73746C756166656420676E",
    INIT_0c => x"00000000000000000000000000000000000001004E0008000050183A000803FF",
    INIT_0d => x"BD0FC625002610B5DF7DE2E7FDA2E7FD1B00CC00000000000000000000000000",
    INIT_0e => x"FD05EC85303D07C64444440235A2E7FD05EC85303D07C65EFF8E0F840234F1F3",
    INIT_0f => x"9DDF8E0F26B5DF7D80A7038680A7FF8680A7018680A700869DDF8EAAF617E2E7",
    INIT_10 => x"470927100FF917E60A17032790F817152A80E7B6F62614C15C80A7F1F3BD10C6",
    INIT_11 => x"B1F3BD21E8BD891FB1F3BD21E8BDF9F2BDA8F28EF9F2BD7EF28E410916F20717",
    INIT_12 => x"F28ECE20F9F2BDADF28EF126FF8184A60230946E022681AC1061F48E021F891E",
    INIT_13 => x"0D0A8ADF9F6E88DF9F6E86DF9F6E84DF9F6E82DF9F6E39A4F07E501A00F3BDC2",
    INIT_14 => x"32206C6C61626D75522E412E442020302E35207265562039306E6F4D202B2B2B",
    INIT_15 => x"21646E616D6D6F63206E776F6E6B6E55200707043E3D0D0A042B2B2B20353030",
    INIT_16 => x"215450555245544E492044455443455058454E55070707070707070707070420",
    INIT_17 => x"39F726048180A623E8BD9035058DEAF28E1034040D0A04212121212121212121",
    INIT_18 => x"10363496356A8D92DF8E92DFBF16349635788D91DF8E91DFB7163439F58DEB8D",
    INIT_19 => x"484848218D043439011F891E058D891F098DB635F3261F30FB263F313DE2048E",
    INIT_1a => x"E8BD23E87E078BCAF423103981308B0F84444444448435E0AB0434198D891F48",
    INIT_1b => x"8D84A6E12023E8BD0886390780032E1681072B11810A2F09810F2B30804E8D21",
    INIT_1c => x"98DF7948489BDFB84848489BDFB608C6043423E87E2086F48DF68DCA2080A6CA",
    INIT_1d => x"02340434392080022E7A81062D6181843598DFB6E6265A9BDF799ADF7999DF79",
    INIT_1e => x"8BF9205C032B0A805F0434843591DFBB91DFF70FC40435981F3D0AC644444444",
    INIT_1f => x"F917981F9AF91740F917D08600F91796351634843591DFBB91DFF7585858580A",
    INIT_20 => x"1702349635163439F8F817A0F91751F91787F9172DF917D186EDF81792F91738",
    INIT_21 => x"123439D3F8175CF91702F917023564F9170AF917981F6CF91712F917D086D2F8",
    INIT_22 => x"6EC1E7B7C0E7B74F923580E7B7F78480E7B61DF3BD19008E80E7B7088A80E7B6",
    INIT_23 => x"F4554A3FF54F5318F54953DBFE425372F64D467CF74D50D3F7454D01F7554484",
    INIT_24 => x"F9535267FB4F4256F84D5414F652448DF54B42CCF5504364F55052F7F4464AD0",
    INIT_25 => x"706D754A0808FFFAFC504C37FC534C4AFE434D73FD434410FA465289F9535714",
    INIT_26 => x"754A080858F47E2EF3BDF9F2BDBAF48E04207461206D6172676F7270206F7420",
    INIT_27 => x"03CD8EF9F2BDDCF48E042E7472617473206D7261772078656C66206F7420706D",
    INIT_28 => x"F3BDF9F2BD03F58E04206F742074726F70207475706E6920746553080858F47E",
    INIT_29 => x"8E04206F742074726F702074757074756F2074655308082CF27E8CDFB703845E",
    INIT_2a => x"7266206D6172676F7270206E755208082CF27E8DDFB703845EF3BDF9F2BD29F5",
    INIT_2b => x"72622074655308083B80DFFE10E4A7FF866AAF2EF3BDF9F2BD50F58E04206D6F",
    INIT_2c => x"7E84A73F86CDDFB784A62EF3BDF9F2BD78F58E0420746120746E696F706B6165",
    INIT_2d => x"662065756E69746E6F4308081AF67E84A7CDDFB66AAF1F306AAE80DFFF102CF2",
    INIT_2e => x"432079616C70736944080873F57EF9F2BDB4F58E042E2E2E2E495753206D6F72",
    INIT_2f => x"202020582050442042202041202043430D0A042E737265747369676572205550",
    INIT_30 => x"F9F2BDEEF58EF9F2BDD5F58E040D0A5320202020435020202055202020205920",
    INIT_31 => x"85F3BD80DF8E85F3BD85F3BD85F3BD85F3BD87F3BD87F3BD87F3BD87F3BD411F",
    INIT_32 => x"6620746E6174736E6F6320687469772079726F6D656D206C6C694608082CF27E",
    INIT_33 => x"65F68E121F2EF3BDF9F2BD43F68E042065756C61762004206F742004206D6F72",
    INIT_34 => x"4808082CF27E1035F926E4AC10A0A739F3BDF9F2BD6AF68E10342EF3BDF9F2BD",
    INIT_35 => x"202030202020202004206D6F72662079726F6D656D20666F20706D7564207865",
    INIT_36 => x"4220204120203920203820202037202036202035202034202033202032202031",
    INIT_37 => x"4645444342413938373635343332313020202020462020452020442020432020",
    INIT_38 => x"F2BD103500F3BDB8F68E1034EDF2BD10008E10EDF2BD2EF3BDF9F2BD9DF68E04",
    INIT_39 => x"A6103010C689F3BD89F3BDF12089F3BDF62608C109275A87F3BD10C611F3BDED",
    INIT_3a => x"2D81AF270D8121E8BDC7263F31EC2002275A23E8BD2E86022D7F81042D208180",
    INIT_3b => x"BD6AF78E042074612079726F6D656D20656B6F500808A32000FE8930C8FA2610",
    INIT_3c => x"78652079726F6D654D08082CF27EA4A739F3BDF9F2BD6AF68E121F2EF3BDF9F2",
    INIT_3d => x"6172206F4E2020070704206D6F726620796669646F6D20646E6120656E696D61",
    INIT_3e => x"BDEDF2BD2EF3BDF9F2BD95F78E0421737365726464612074616874207461206D",
    INIT_3f => x"A11FA739F3BD32FA26102081E8270D81EC201E3004262D8121E8BD87F3BD11F3"


	 )

   port map (
      DO => rdata1,                -- 8-bit Data Output
      DOP => dp1,                  -- 1-bit parity Output
      ADDR => addr(10 downto 0),   -- 11-bit Address Input
      CLK => clk,                  -- Clock
      DI => wdata,                 -- 8-bit Data Input
      DIP => dp1,                  -- 1-bit parity Input
      EN => cs1,                   -- RAM Enable Input
      SSR => rst,                  -- Synchronous Set/Reset Input
      WE => we                     -- Write Enable Input
   );
   -- End of RAMB16_S9_inst instantiation
 
   RAM_2 : RAMB16_S9	-- $F800 - $FFFF
   generic map (
      INIT => X"000", --  Value of output RAM registers at startup
      SRVAL => X"000", --  Ouput value upon SSR assertion
      WRITE_MODE => "WRITE_FIRST", --  WRITE_FIRST, READ_FIRST or NO_CHANGE
    INIT_00 => x"04206D6F72662079726F6D656D207473655408082CF27EF9F2BDB7F78ED9271F",
    INIT_01 => x"74206465676E61686304206E6F697461636F6C20746120726F7272450D0A0707",
    INIT_02 => x"1F2EF3BDF9F2BD0CF88E04206874697720776F6E20676E69747365542004206F",
    INIT_03 => x"E7211F7DF3BD91DF8E91DFF7F9F2BD43F88E5F92DFBF2EF3BDF9F2BD65F68E12",
    INIT_04 => x"8E2CF27ED820121F23E8BD23E8BD08860C275CF22692DFBC1021311A26A4E1A4",
    INIT_05 => x"F88E87F3BD91DF8E91DFF789F3BD89F3BD85F3BD92DF8E92DFBF10F9F2BD20F8",
    INIT_06 => x"636573206D6F726620646165520808CB2087F3BD91DF8E91DFB7A4A6F9F2BD37",
    INIT_07 => x"0D0420726F746365732004206B636172742004206576697264206E6F20726F74",
    INIT_08 => x"8EDFB75EF3BDF9F2BDD1F88E04203D2065646F6320726F72726520434446070A",
    INIT_09 => x"F68E90DFB739F3BDF9F2BDF6F88E8FDFB739F3BDF9F2BDEEF88E99ECBD8BDF8E",
    INIT_0a => x"91DF8E91DFF7F9F2BDFFF88ED8F8271084ECBD90DFF68FDFB62EF3BDF9F2BD65",
    INIT_0b => x"6576697264206E6F20726F74636573206F7420657469725708082CF27E87F3BD",
    INIT_0c => x"F2BDEEF88E99ECBD8BDF8E8EDFB75EF3BDF9F2BD66F98E04206D6F7266200420",
    INIT_0d => x"F68FDFB62EF3BDF9F2BD82F98E90DFB739F3BDF9F2BDF6F88E8FDFB739F3BDF9",
    INIT_0e => x"726F4608082CF27E87F3BD91DF8E91DFF7F9F2BDFFF88E63F8271088ECBD90DF",
    INIT_0f => x"6F6E206B7369646D615207040D0A202E2E2E6B7369644D415220676E6974616D",
    INIT_10 => x"A65F9DDF8EF9F2BDDBF98E17F816038D040D0A202164657461636F6C6C612074",
    INIT_11 => x"A75F4F80DE8E99ECBD8BDF8E8EDFF73900F3BDF5F98EF52604C15C0C27018180",
    INIT_12 => x"0186846C042625814C90DFB684A78FDFB680DE8E90DFB701868FDF7FFB265A80",
    INIT_13 => x"8FDFB68FDF7C90DFB70186D726258190DFB690DF7C88ECBD90DFF68FDFB601A7",
    INIT_14 => x"4F80DE8E88ECBD24C64F86016F846F80DE8E84ECBD24C64F8680DE8EC8265081",
    INIT_15 => x"846F80DE8E84ECBD03C64F80DE8E88ECBD24C64F016F846F80DE8E84ECBD24C6",
    INIT_16 => x"1B88ED0100CC1688ED204BCC1488ED5349CC1288ED444DCC1088ED4152CC016F",
    INIT_17 => x"862488A71F862388A701862188ED1C0BCC2688ED1F88ED244FCC1D88ED0101CC",
    INIT_18 => x"C62488A7BCF3BDF1F3BD04C62388A7BCF3BDF1F3BD05C62126B5DF7D2588A705",
    INIT_19 => x"84A7AA8680DE8E84ECBD01C64F80DE8E88ECBD03C64F2588A7BCF3BDF1F3BD06",
    INIT_1a => x"4C46206C616E7265746E6920676E69746F6F4208083988ECBD01C64F01A75586",
    INIT_1b => x"00DE8EF726FDD38C81EDA1ECCDFB8E10E5D38EF9F2BD4BFB8E042E2E2E2E5845",
    INIT_1c => x"B7BCF3BDF1F3BD05C602CAB739863526B5DF7DF7261EDE8C81EDA1ECE5FB8E10",
    INIT_1d => x"F1F3BD14C600CC8E10CCB7BCF3BDF1F3BD06C60FCCB7BCF3BDF1F3BD04C60ECC",
    INIT_1e => x"E869F22CF269F269F269F2FEFFFEFF69F210E858F47E00CD8EF62621C15C80A7",
    INIT_1f => x"ECEC7ED4EC7ED0EC7ECCEC7E99EC7E90EC7E8CEC7E88EC7E84EC7E21E823E800",
    INIT_20 => x"6420726F6620676E6974696177202C6B7369644D4F522064616F4C0808F0EC7E",
    INIT_21 => x"028E10F9F2BD03FC8E040808080808042020202020202E2E2E64616F6C6E776F",
    INIT_22 => x"D2E7F73FC4101F00FE8930211F1034F8265A80A788FCBD5FC0E7BF1000008E00",
    INIT_23 => x"008E10C42600048C1021311035D3E7B791DFBB484891DFF7545454545454101F",
    INIT_24 => x"354DE8BD04348435E0AB0434068D891F484848480E8D04342CF27EC0E7BF1000",
    INIT_25 => x"69644D4F522064616F4C0808390780E92E1681ED2B11810A2F0981F52B308004",
    INIT_26 => x"4E595320646E756F462020042E4D4F5250206769666E6F63206D6F7266206B73",
    INIT_27 => x"8E2DF516038D040D0A2E2E2E6174616420676E6964616F6C202C64726F772043",
    INIT_28 => x"8E10F9F2BDD5FC8EF9270184F1E7B60CF61764008EF2E7B7F0E7B6F9F2BDB4FC",
    INIT_29 => x"2600048C102131F1265A80A7F0E7B6F9270284F1E7B65FC0E7BF1000008E0002",
    INIT_2a => x"2E73746E65746E6F63204354522079616C707369440D39C0E7BF1000008E10E1",
    INIT_2b => x"FD8E0927B5DF7DF9F2BD4AFD8E0421646E756F6620435452206F4E2020200704",
    INIT_2c => x"8620FEBDF1F3BD01C623E8BD3A8620FEBDF1F3BD02C6EDF2BD2CF27EF9F2BD61",
    INIT_2d => x"BD2F86638DF1F3BD04C623E8BD208623E8BD208620FEBDF1F3BD00C623E8BD3A",
    INIT_2e => x"C6288D06008E08C6EDF2BD4B8DF1F3BD06C623E8BD2F86578DF1F3BD05C623E8",
    INIT_2f => x"8E088D0F008E0D8D02008E128D0B008E178D04008E1C8D01008E218D01008E0E",
    INIT_30 => x"39EDF2BDEB261F30103587F3BD91DF8E103491DFB75CF1F3BD2CF27E038D1000",
    INIT_31 => x"6C6120646E6120656E696D617865204354520D96357DF3BD91DF8E91DFB71634",
    INIT_32 => x"F3BD2CF27EF9F2BD61FD8E0927B5DF7DF9F2BD2DFE8E04206D6F726620726574",
    INIT_33 => x"21E8BD7DF3BD91DF8E91DFB7F1F3BD87F3BD91DF8E91DFF7EDF2BD3FC4891F39",
    INIT_34 => x"530808C6205A92F326102D81CF205C03260D81D6205C1DF4BD39F3BD09262081",
    INIT_35 => x"74617220647561622004206169636120726F6620657461722064756162207465",
    INIT_36 => x"F2BD9DFE8E042E6E776F6E6B20746F6E206574617220647561422004203D2065",
    INIT_37 => x"105F5EFF8E021E891E21E8BD891F21E8BDF9F2BDB7FE8E91DFB701845EF3BDF9",
    INIT_38 => x"E8BD03A623E8BD02A604342CF27EF9F2BDC5FE8EF32696FF8C5C0730112784AC",
    INIT_39 => x"BAF08491DFF70435A2E7BF1010265D91DFF605AE10F1F3BD0FC623E8BD04A623",
    INIT_3a => x"30332CF27E1DF4BD0FC691DFBA0F8491DFF7585858580435E2E7BF10122091DF",
    INIT_3b => x"002030303639460120303038348B022030303432160520303032315814202030",
    INIT_3c => x"000000000000000000FF1B0030303637352900303034383351003030323931A3",
    INIT_3d => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3e => x"F27E69F27E69F27E69F27E69F27E69F27E69F27E69F27E23E87E10E87E00E87E",
    INIT_3f => x"A4F06AF2A2F56EF272F276F27AF2A4F069F27E69F27E69F27E69F27E69F27E69"




	 )

   port map (
      DO => rdata2,                -- 8-bit Data Output
      DOP => dp2,                  -- 1-bit parity Output
      ADDR => addr(10 downto 0),   -- 11-bit Address Input
      CLK => clk,                  -- Clock
      DI => wdata,                 -- 8-bit Data Input
      DIP => dp2,                  -- 1-bit parity Input
      EN => cs2,                   -- RAM Enable Input
      SSR => rst,                  -- Synchronous Set/Reset Input
      WE => we                     -- Write Enable Input
   );
   -- End of RAMB16_S9_inst instantiation


   -- Decode high order address bits to select block, mux data outputs
   decode_and_data_mux : process (addr(12 downto 11),
                                  cs0, cs1, cs2 )  
   begin
   	we <= not rw;
   	case addr(12 downto 11) is
	
		-- $F800 - $FFFF
		when "11" => 
		   rdata <= rdata2;
		   cs2 <= cs; 
		   cs1 <= '0';
		   cs0 <= '0';
 
		-- $F000 - $F7FF
		when "10" => 
		   rdata <= rdata1;
		   cs2 <= '0'; 
		   cs1 <= cs;
		   cs0 <= '0';

		-- $E800 - EFFF
		when "01" => 
		   rdata <= rdata0; 
		   cs2 <= '0'; 
		   cs1 <= '0';
		   cs0 <= cs;

		-- $E000 - E7FF  (external to this ROM - screen buffer and IO space)
		when others => 
		   rdata <= rdata0;   -- data is 'don't care' at this point
		   cs2 <= '0'; 
		   cs1 <= '0';
		   cs0 <= '0';

	end case;
			      
   end process;

end architecture;
