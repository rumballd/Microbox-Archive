----------------------------------------------------------------
--
-- Character generator ROM - definitions from MB2 'pretty' char set
--
-- 7 pixels x 11 rows x 128 characters.	
-- organised as 8x16, top row and bottom four rows blank.
-- (using new Xilinx component definitions)
----------------------------------------------------------------

library IEEE, UNISIM;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use UNISIM.vcomponents.all;

entity char_rom is
    Port (
     clk   : in  std_logic;
	rst   : in  std_logic;
	cs    : in  std_logic;
	rw    : in  std_logic;
     addr  : in  std_logic_vector (10 downto 0);
     rdata : out std_logic_vector (7 downto 0);
     wdata : in  std_logic_vector (7 downto 0)
    );

end char_rom;

architecture rtl of char_rom is

   signal dp : std_logic_vector(0 downto 0);	-- loop parity bit output to input

begin
   
   RAM_0 : RAMB16_S9
   generic map (
      INIT => X"000", --  Value of output RAM registers at startup
      SRVAL => X"000", --  Ouput value upon SSR assertion
      WRITE_MODE => "WRITE_FIRST", --  WRITE_FIRST, READ_FIRST or NO_CHANGE
    INIT_00 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_01 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_02 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_03 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_04 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_05 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_06 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_07 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_08 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_09 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0a => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0b => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0c => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0d => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0e => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0f => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_10 => x"0000000000000008080008080808080000000000000000000000000000000000",
    INIT_11 => x"0000000000001414147F147F1414140000000000000000000000000024242400",
    INIT_12 => x"00000000000002452210080422512000000000000000087E09093E48483F0800",
    INIT_13 => x"000000000000000000000010080C0C0000000000000039464629102844443800",
    INIT_14 => x"0000000000001008040404040408100000000000000004081010101010080400",
    INIT_15 => x"000000000000000808087F08080800000000000000000008492A7F2A49080000",
    INIT_16 => x"000000000000000000003E000000000000000000201018180000000000000000",
    INIT_17 => x"0000000000000040201008040201000000000000000018180000000000000000",
    INIT_18 => x"0000000000003E0808080808281808000000000000003E416151494543413E00",
    INIT_19 => x"0000000000003E4101011E0101413E000000000000007F4040201C0201413E00",
    INIT_1a => x"0000000000003C420101027C40407F0000000000000002027F4222120A060200",
    INIT_1b => x"00000000000010101010080402417F000000000000003E4141417E4040201E00",
    INIT_1c => x"0000000000003C0201013F4141413E000000000000003E4141413E4141413E00",
    INIT_1d => x"0000000020101818000018180000000000000000000018180000181800000000",
    INIT_1e => x"0000000000000000003E003E0000000000000000000004081020402010080400",
    INIT_1f => x"00000000000008000808060121211E0000000000000010080402010204081000",
    INIT_20 => x"0000000000004141417F414141221C000000000000001E20405E55554D211E00",
    INIT_21 => x"0000000000001E214040404040211E000000000000007E2121213E2121217E00",
    INIT_22 => x"0000000000007F404040784040407F000000000000007C424141414141427C00",
    INIT_23 => x"0000000000001E21414F404040211E0000000000000040404040784040407F00",
    INIT_24 => x"0000000000003E080808080808083E00000000000000414141417F4141414100",
    INIT_25 => x"0000000000004142446850484442410000000000000038440404040404041F00",
    INIT_26 => x"000000000000414141414949556341000000000000007F404040404040404000",
    INIT_27 => x"0000000000001C224141414141221C0000000000000041414143454951614100",
    INIT_28 => x"0000000000001D224549414141221C00000000000000404040407E4141417E00",
    INIT_29 => x"0000000000003E4101013E4040413E00000000000000414244487E4141417E00",
    INIT_2a => x"0000000000003E41414141414141410000000000000008080808080808087F00",
    INIT_2b => x"0000000000004163554949414141410000000000000008081414222241414100",
    INIT_2c => x"0000000000000808080808142241410000000000000041412214081422414100",
    INIT_2d => x"0000000000003E202020202020203E000000000000007F402010080402017F00",
    INIT_2e => x"0000000000003E020202020202023E0000000000000000010204081020400000",
    INIT_2f => x"0000000000003E0000000000000000000000000000000808080808492A1C0800",
    INIT_30 => x"0000000000003D42423E023C0000000000000000000000000000000408181800",
    INIT_31 => x"0000000000003C424040423C000000000000000000005C624242625C40404000",
    INIT_32 => x"0000000000003C40407E423C000000000000000000003A464242463A02020200",
    INIT_33 => x"000000003C42023A4642463A00000000000000000000101010107C1010120C00",
    INIT_34 => x"0000000000001C08080808180008000000000000000042424242625C40404000",
    INIT_35 => x"00000000000042446850484440404000000000001C2202020202020600020000",
    INIT_36 => x"000000000000494949494976000000000000000000001C080808080808081800",
    INIT_37 => x"0000000000003E414141413E0000000000000000000042424242625C00000000",
    INIT_38 => x"000000000302023A4642463A00000000000000004040405C6242625C00000000",
    INIT_39 => x"0000000000003C420C30423C0000000000000000000040404040625C00000000",
    INIT_3a => x"0000000000003A4642424242000000000000000000000C121010107C10100000",
    INIT_3b => x"0000000000003649494949410000000000000000000008142241414100000000",
    INIT_3c => x"000000003C42023A464242420000000000000000000042241818244200000000",
    INIT_3d => x"0000000000000C101010201010100C000000000000007E201008047E00000000",
    INIT_3e => x"0000000000001804040402040404180000000000000000000808080008080800",
    INIT_3f => x"0000000000002A552A552A552A552A0000000000000000000000000006493000"

	 )

   port map (
      DO => rdata,                 -- 8-bit Data Output
      DOP => dp,                   -- 1-bit parity Output
      ADDR => addr(10 downto 0),   -- 11-bit Address Input
      CLK => clk,                  -- Clock
      DI => wdata,                 -- 8-bit Data Input
      DIP => dp,                   -- 1-bit parity Input
      EN => cs,                    -- RAM Enable Input
      SSR => rst,                  -- Synchronous Set/Reset Input
      WE => not rw                 -- Write Enable Input
   );
   -- End of RAMB16_S9_inst instantiation

end architecture rtl;

